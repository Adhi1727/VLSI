module seq_dec(
input clk,rst,x,
output z
);
parameter s0 = 3'b000;
parameter s1 = 3'b001;
parameter s2 = 3'b010;
parameter s3 = 3'b011;
parameter s4 = 3'b100;

reg [2:0] state,next_state;

always @(posedge clk ) begin
	if (!rst) begin 
		state <= s0;
	end
	else
		state <= next_state;
end

	always @(state or x) begin
		case(state) 
	        s0:begin
		if(x==0) next_state = s1;
		else next_state = s3;
		end

		s1:begin
		if(x==0) next_state = s2;
		else next_state = s3;
		end

		s2:begin
		if(x==0) next_state = s2;
		else next_state = s3;
		end

		s3:begin
		if(x==1) next_state = s4;
		else next_state = s1;
		end

		s4:begin
		if(x==1) next_state = s4;
		else next_state = s1;
		end
		default: next_state = s0;
		endcase
		
	end
	assign z = ( ((state==s4)&&(x==1)) || ((state==s2)&&(x==0)) )? 1:0;
endmodule
