module and_opr(
input a,b,
output y
);

	assign y = a&b;
endmodule
