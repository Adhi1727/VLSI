module not_sys(
    input a,
    output y
);
    assign y = ~a;
endmodule

